/*###########################################################*/
/*                 Clock and reset assign                    */
/*                                                           */
/*###########################################################*/
 wire axi_fabric_clk;
 wire axi_fabric_rst_n;
 
 assign axi_fabric_clk = clk;
 assign axi_fabric_rst_n = rstn;
 
 
/*###########################################################*/
/*                 axi_fabric_top_wrapper interface                   */
/*                       (Vtool)                             */
/*###########################################################*/
   axi_fabric_top_wrapper
    #(
       .SLAVE_N(),
       .MASTER_N(),
       .ADDR_WIDTH(),
       .DATA_WIDTH(),
       .S_ID_WIDTH(),
       .M_ID_WIDTH(),
       .STRB_WIDTH(),
       .AW_USER_WIDTH(),
       .W_USER_WIDTH(),
       .B_USER_WIDTH(),
       .AR_USER_WIDTH(),
       .R_USER_WIDTH(),
       .ARBITER_TYPE(),
       .MAX_TRANS(),
       .S_AR_CHANNEL_REG(),
       .M_AR_CHANNEL_REG(),
       .S_R_CHANNEL_REG(),
       .M_R_CHANNEL_REG(),
       .S_AW_CHANNEL_REG(),
       .M_AW_CHANNEL_REG(),
       .S_W_CHANNEL_REG(),
       .M_W_CHANNEL_REG(),
       .S_WR_CHANNEL_REG(),
       .M_WR_CHANNEL_REG()
   )
   axi_fabric_top_wrapper_inst (
        .clk(clk),
        .rst_n(rst_n),
        .s00_axi_awid(s00_axi_awid),
        .s00_axi_awaddr(s00_axi_awaddr),
        .s00_axi_awlen(s00_axi_awlen),
        .s00_axi_awsize(s00_axi_awsize),
        .s00_axi_awburst(s00_axi_awburst),
        .s00_axi_awlock(s00_axi_awlock),
        .s00_axi_awcache(s00_axi_awcache),
        .s00_axi_awprot(s00_axi_awprot),
        .s00_axi_awqos(s00_axi_awqos),
        .s00_axi_awuser(s00_axi_awuser),
        .s00_axi_awvalid(s00_axi_awvalid),
        .s00_axi_awready(s00_axi_awready),
        .s00_axi_wdata(s00_axi_wdata),
        .s00_axi_wstrb(s00_axi_wstrb),
        .s00_axi_wuser(s00_axi_wuser),
        .s00_axi_wvalid(s00_axi_wvalid),
        .s00_axi_wready(s00_axi_wready),
        .s00_axi_wlast(s00_axi_wlast),
        .s00_axi_bid(s00_axi_bid),
        .s00_axi_buser(s00_axi_buser),
        .s00_axi_bresp(s00_axi_bresp),
        .s00_axi_bvalid(s00_axi_bvalid),
        .s00_axi_bready(s00_axi_bready),
        .s00_axi_arid(s00_axi_arid),
        .s00_axi_araddr(s00_axi_araddr),
        .s00_axi_aruser(s00_axi_aruser),
        .s00_axi_arlen(s00_axi_arlen),
        .s00_axi_arsize(s00_axi_arsize),
        .s00_axi_arburst(s00_axi_arburst),
        .s00_axi_arlock(s00_axi_arlock),
        .s00_axi_arcache(s00_axi_arcache),
        .s00_axi_arprot(s00_axi_arprot),
        .s00_axi_arqos(s00_axi_arqos),
        .s00_axi_arvalid(s00_axi_arvalid),
        .s00_axi_arready(s00_axi_arready),
        .s00_axi_rdata(s00_axi_rdata),
        .s00_axi_rid(s00_axi_rid),
        .s00_axi_rresp(s00_axi_rresp),
        .s00_axi_rlast(s00_axi_rlast),
        .s00_axi_rvalid(s00_axi_rvalid),
        .s00_axi_ruser(s00_axi_ruser),
        .s00_axi_rready(s00_axi_rready),
        .s01_axi_awid(s01_axi_awid),
        .s01_axi_awaddr(s01_axi_awaddr),
        .s01_axi_awuser(s01_axi_awuser),
        .s01_axi_awlen(s01_axi_awlen),
        .s01_axi_awsize(s01_axi_awsize),
        .s01_axi_awburst(s01_axi_awburst),
        .s01_axi_awlock(s01_axi_awlock),
        .s01_axi_awcache(s01_axi_awcache),
        .s01_axi_awprot(s01_axi_awprot),
        .s01_axi_awqos(s01_axi_awqos),
        .s01_axi_awvalid(s01_axi_awvalid),
        .s01_axi_awready(s01_axi_awready),
        .s01_axi_wdata(s01_axi_wdata),
        .s01_axi_wuser(s01_axi_wuser),
        .s01_axi_wstrb(s01_axi_wstrb),
        .s01_axi_wvalid(s01_axi_wvalid),
        .s01_axi_wready(s01_axi_wready),
        .s01_axi_wlast(s01_axi_wlast),
        .s01_axi_bid(s01_axi_bid),
        .s01_axi_buser(s01_axi_buser),
        .s01_axi_bresp(s01_axi_bresp),
        .s01_axi_bvalid(s01_axi_bvalid),
        .s01_axi_bready(s01_axi_bready),
        .s01_axi_arid(s01_axi_arid),
        .s01_axi_araddr(s01_axi_araddr),
        .s01_axi_aruser(s01_axi_aruser),
        .s01_axi_arlen(s01_axi_arlen),
        .s01_axi_arsize(s01_axi_arsize),
        .s01_axi_arburst(s01_axi_arburst),
        .s01_axi_arlock(s01_axi_arlock),
        .s01_axi_arcache(s01_axi_arcache),
        .s01_axi_arprot(s01_axi_arprot),
        .s01_axi_arqos(s01_axi_arqos),
        .s01_axi_arvalid(s01_axi_arvalid),
        .s01_axi_arready(s01_axi_arready),
        .s01_axi_rdata(s01_axi_rdata),
        .s01_axi_rid(s01_axi_rid),
        .s01_axi_rresp(s01_axi_rresp),
        .s01_axi_rlast(s01_axi_rlast),
        .s01_axi_rvalid(s01_axi_rvalid),
        .s01_axi_ruser(s01_axi_ruser),
        .s01_axi_rready(s01_axi_rready),
        .s02_axi_awid(s02_axi_awid),
        .s02_axi_awaddr(s02_axi_awaddr),
        .s02_axi_awuser(s02_axi_awuser),
        .s02_axi_awlen(s02_axi_awlen),
        .s02_axi_awsize(s02_axi_awsize),
        .s02_axi_awburst(s02_axi_awburst),
        .s02_axi_awlock(s02_axi_awlock),
        .s02_axi_awcache(s02_axi_awcache),
        .s02_axi_awprot(s02_axi_awprot),
        .s02_axi_awqos(s02_axi_awqos),
        .s02_axi_awvalid(s02_axi_awvalid),
        .s02_axi_awready(s02_axi_awready),
        .s02_axi_wdata(s02_axi_wdata),
        .s02_axi_wuser(s02_axi_wuser),
        .s02_axi_wstrb(s02_axi_wstrb),
        .s02_axi_wvalid(s02_axi_wvalid),
        .s02_axi_wready(s02_axi_wready),
        .s02_axi_wlast(s02_axi_wlast),
        .s02_axi_bid(s02_axi_bid),
        .s02_axi_buser(s02_axi_buser),
        .s02_axi_bresp(s02_axi_bresp),
        .s02_axi_bvalid(s02_axi_bvalid),
        .s02_axi_bready(s02_axi_bready),
        .s02_axi_arid(s02_axi_arid),
        .s02_axi_araddr(s02_axi_araddr),
        .s02_axi_aruser(s02_axi_aruser),
        .s02_axi_arlen(s02_axi_arlen),
        .s02_axi_arsize(s02_axi_arsize),
        .s02_axi_arburst(s02_axi_arburst),
        .s02_axi_arlock(s02_axi_arlock),
        .s02_axi_arcache(s02_axi_arcache),
        .s02_axi_arprot(s02_axi_arprot),
        .s02_axi_arqos(s02_axi_arqos),
        .s02_axi_arvalid(s02_axi_arvalid),
        .s02_axi_arready(s02_axi_arready),
        .s02_axi_rdata(s02_axi_rdata),
        .s02_axi_rid(s02_axi_rid),
        .s02_axi_rresp(s02_axi_rresp),
        .s02_axi_rlast(s02_axi_rlast),
        .s02_axi_rvalid(s02_axi_rvalid),
        .s02_axi_ruser(s02_axi_ruser),
        .s02_axi_rready(s02_axi_rready),
        .m00_axi_awid(m00_axi_awid),
        .m00_axi_awaddr(m00_axi_awaddr),
        .m00_axi_awlen(m00_axi_awlen),
        .m00_axi_awsize(m00_axi_awsize),
        .m00_axi_awburst(m00_axi_awburst),
        .m00_axi_awlock(m00_axi_awlock),
        .m00_axi_awcache(m00_axi_awcache),
        .m00_axi_awprot(m00_axi_awprot),
        .m00_axi_awregion(m00_axi_awregion),
        .m00_axi_awqos(m00_axi_awqos),
        .m00_axi_awuser(m00_axi_awuser),
        .m00_axi_awvalid(m00_axi_awvalid),
        .m00_axi_awready(m00_axi_awready),
        .m00_axi_wdata(m00_axi_wdata),
        .m00_axi_wstrb(m00_axi_wstrb),
        .m00_axi_wuser(m00_axi_wuser),
        .m00_axi_wvalid(m00_axi_wvalid),
        .m00_axi_wready(m00_axi_wready),
        .m00_axi_wlast(m00_axi_wlast),
        .m00_axi_bid(m00_axi_bid),
        .m00_axi_buser(m00_axi_buser),
        .m00_axi_bresp(m00_axi_bresp),
        .m00_axi_bvalid(m00_axi_bvalid),
        .m00_axi_bready(m00_axi_bready),
        .m00_axi_araddr(m00_axi_araddr),
        .m00_axi_arid(m00_axi_arid),
        .m00_axi_arlen(m00_axi_arlen),
        .m00_axi_arsize(m00_axi_arsize),
        .m00_axi_arburst(m00_axi_arburst),
        .m00_axi_arlock(m00_axi_arlock),
        .m00_axi_arcache(m00_axi_arcache),
        .m00_axi_arprot(m00_axi_arprot),
        .m00_axi_arregion(m00_axi_arregion),
        .m00_axi_arqos(m00_axi_arqos),
        .m00_axi_aruser(m00_axi_aruser),
        .m00_axi_arvalid(m00_axi_arvalid),
        .m00_axi_arready(m00_axi_arready),
        .m00_axi_rdata(m00_axi_rdata),
        .m00_axi_rid(m00_axi_rid),
        .m00_axi_rresp(m00_axi_rresp),
        .m00_axi_rlast(m00_axi_rlast),
        .m00_axi_rvalid(m00_axi_rvalid),
        .m00_axi_ruser(m00_axi_ruser),
        .m00_axi_rready(m00_axi_rready),
        .m01_axi_awid(m01_axi_awid),
        .m01_axi_awaddr(m01_axi_awaddr),
        .m01_axi_awlen(m01_axi_awlen),
        .m01_axi_awsize(m01_axi_awsize),
        .m01_axi_awburst(m01_axi_awburst),
        .m01_axi_awlock(m01_axi_awlock),
        .m01_axi_awcache(m01_axi_awcache),
        .m01_axi_awprot(m01_axi_awprot),
        .m01_axi_awregion(m01_axi_awregion),
        .m01_axi_awqos(m01_axi_awqos),
        .m01_axi_awuser(m01_axi_awuser),
        .m01_axi_awvalid(m01_axi_awvalid),
        .m01_axi_awready(m01_axi_awready),
        .m01_axi_wdata(m01_axi_wdata),
        .m01_axi_wstrb(m01_axi_wstrb),
        .m01_axi_wuser(m01_axi_wuser),
        .m01_axi_wvalid(m01_axi_wvalid),
        .m01_axi_wready(m01_axi_wready),
        .m01_axi_wlast(m01_axi_wlast),
        .m01_axi_bid(m01_axi_bid),
        .m01_axi_buser(m01_axi_buser),
        .m01_axi_bresp(m01_axi_bresp),
        .m01_axi_bvalid(m01_axi_bvalid),
        .m01_axi_bready(m01_axi_bready),
        .m01_axi_araddr(m01_axi_araddr),
        .m01_axi_arid(m01_axi_arid),
        .m01_axi_arlen(m01_axi_arlen),
        .m01_axi_arsize(m01_axi_arsize),
        .m01_axi_arburst(m01_axi_arburst),
        .m01_axi_arlock(m01_axi_arlock),
        .m01_axi_arcache(m01_axi_arcache),
        .m01_axi_arprot(m01_axi_arprot),
        .m01_axi_arregion(m01_axi_arregion),
        .m01_axi_arqos(m01_axi_arqos),
        .m01_axi_aruser(m01_axi_aruser),
        .m01_axi_arvalid(m01_axi_arvalid),
        .m01_axi_arready(m01_axi_arready),
        .m01_axi_rdata(m01_axi_rdata),
        .m01_axi_rid(m01_axi_rid),
        .m01_axi_rresp(m01_axi_rresp),
        .m01_axi_rlast(m01_axi_rlast),
        .m01_axi_rvalid(m01_axi_rvalid),
        .m01_axi_ruser(m01_axi_ruser),
        .m01_axi_rready(m01_axi_rready),
        .m02_axi_awid(m02_axi_awid),
        .m02_axi_awaddr(m02_axi_awaddr),
        .m02_axi_awlen(m02_axi_awlen),
        .m02_axi_awsize(m02_axi_awsize),
        .m02_axi_awburst(m02_axi_awburst),
        .m02_axi_awlock(m02_axi_awlock),
        .m02_axi_awcache(m02_axi_awcache),
        .m02_axi_awprot(m02_axi_awprot),
        .m02_axi_awregion(m02_axi_awregion),
        .m02_axi_awqos(m02_axi_awqos),
        .m02_axi_awuser(m02_axi_awuser),
        .m02_axi_awvalid(m02_axi_awvalid),
        .m02_axi_awready(m02_axi_awready),
        .m02_axi_wdata(m02_axi_wdata),
        .m02_axi_wstrb(m02_axi_wstrb),
        .m02_axi_wuser(m02_axi_wuser),
        .m02_axi_wvalid(m02_axi_wvalid),
        .m02_axi_wready(m02_axi_wready),
        .m02_axi_wlast(m02_axi_wlast),
        .m02_axi_bid(m02_axi_bid),
        .m02_axi_buser(m02_axi_buser),
        .m02_axi_bresp(m02_axi_bresp),
        .m02_axi_bvalid(m02_axi_bvalid),
        .m02_axi_bready(m02_axi_bready),
        .m02_axi_araddr(m02_axi_araddr),
        .m02_axi_arid(m02_axi_arid),
        .m02_axi_arlen(m02_axi_arlen),
        .m02_axi_arsize(m02_axi_arsize),
        .m02_axi_arburst(m02_axi_arburst),
        .m02_axi_arlock(m02_axi_arlock),
        .m02_axi_arcache(m02_axi_arcache),
        .m02_axi_arprot(m02_axi_arprot),
        .m02_axi_arregion(m02_axi_arregion),
        .m02_axi_arqos(m02_axi_arqos),
        .m02_axi_aruser(m02_axi_aruser),
        .m02_axi_arvalid(m02_axi_arvalid),
        .m02_axi_arready(m02_axi_arready),
        .m02_axi_rdata(m02_axi_rdata),
        .m02_axi_rid(m02_axi_rid),
        .m02_axi_rresp(m02_axi_rresp),
        .m02_axi_rlast(m02_axi_rlast),
        .m02_axi_rvalid(m02_axi_rvalid),
        .m02_axi_ruser(m02_axi_ruser),
        .m02_axi_rready(m02_axi_rready),
        .m03_axi_awid(m03_axi_awid),
        .m03_axi_awaddr(m03_axi_awaddr),
        .m03_axi_awlen(m03_axi_awlen),
        .m03_axi_awsize(m03_axi_awsize),
        .m03_axi_awburst(m03_axi_awburst),
        .m03_axi_awlock(m03_axi_awlock),
        .m03_axi_awcache(m03_axi_awcache),
        .m03_axi_awprot(m03_axi_awprot),
        .m03_axi_awregion(m03_axi_awregion),
        .m03_axi_awqos(m03_axi_awqos),
        .m03_axi_awuser(m03_axi_awuser),
        .m03_axi_awvalid(m03_axi_awvalid),
        .m03_axi_awready(m03_axi_awready),
        .m03_axi_wdata(m03_axi_wdata),
        .m03_axi_wstrb(m03_axi_wstrb),
        .m03_axi_wuser(m03_axi_wuser),
        .m03_axi_wvalid(m03_axi_wvalid),
        .m03_axi_wready(m03_axi_wready),
        .m03_axi_wlast(m03_axi_wlast),
        .m03_axi_bid(m03_axi_bid),
        .m03_axi_buser(m03_axi_buser),
        .m03_axi_bresp(m03_axi_bresp),
        .m03_axi_bvalid(m03_axi_bvalid),
        .m03_axi_bready(m03_axi_bready),
        .m03_axi_araddr(m03_axi_araddr),
        .m03_axi_arid(m03_axi_arid),
        .m03_axi_arlen(m03_axi_arlen),
        .m03_axi_arsize(m03_axi_arsize),
        .m03_axi_arburst(m03_axi_arburst),
        .m03_axi_arlock(m03_axi_arlock),
        .m03_axi_arcache(m03_axi_arcache),
        .m03_axi_arprot(m03_axi_arprot),
        .m03_axi_arregion(m03_axi_arregion),
        .m03_axi_arqos(m03_axi_arqos),
        .m03_axi_aruser(m03_axi_aruser),
        .m03_axi_arvalid(m03_axi_arvalid),
        .m03_axi_arready(m03_axi_arready),
        .m03_axi_rdata(m03_axi_rdata),
        .m03_axi_rid(m03_axi_rid),
        .m03_axi_rresp(m03_axi_rresp),
        .m03_axi_rlast(m03_axi_rlast),
        .m03_axi_rvalid(m03_axi_rvalid),
        .m03_axi_ruser(m03_axi_ruser),
        .m03_axi_rready(m03_axi_rready)
    );

